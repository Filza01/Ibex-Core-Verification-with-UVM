interface dut_intf (input clk);
    bit fetch_enable_i;   // from CPU control signals
    bit reset;
endinterface